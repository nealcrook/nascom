//
module sn74ls161
  (//Out
   output p14,
   output p13,
   output p12,
   output p11,
   // In
   input p1,
   input p2,
   input p7,
   input p9,
   input p10
   );
    initial $display("%m not yet modelled!!");
endmodule // sn74ls161
