//
module x2102an
  (
   output dout,

   input  din,
   input  [9:0] a,
   input  cs_n,
   input  r_nw
   );

    // TODO TEMP
    assign dout = 1'b0;

endmodule // x2102an

