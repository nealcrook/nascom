//
module sn74ls74
  (// Out
   output p9_q,
   output p8_qn,
   // TODO other pair

   // In
   input p11_clk,
   input p12_d,
   input p13_r_n,
   input p10_s_n
   );
    initial $display("%m not yet modelled!!");
endmodule // sn74ls74
