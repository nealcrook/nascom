//
module sn74ls13
  (
   );
    initial $display("%m not yet modelled!!");
endmodule // sn74ls13
