//
module dp8304
  (
   );
    initial $display("%m not yet modelled!!");
endmodule // dp8304

