//
module sn74ls193
  (
   );
    initial $display("%m not yet modelled!!");
endmodule // sn74ls193
