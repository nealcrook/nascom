//
module sn74ls161
  (
   );
    initial $display("%m not yet modelled!!");
endmodule // sn74ls161
