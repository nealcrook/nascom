//
module sn74ls193
  (// Output
   output p13,
   output p12,
   output p7,
   output p6,
   output p2,
   output p3,
   // In
   input  p4,
   input  p1,
   input  p5,
   input  p9,
   input  p10,
   input  p11,
   input  p15,
   input  p14
   );
    initial $display("%m not yet modelled!!");
endmodule // sn74ls193
