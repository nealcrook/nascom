//
module sn74ls74
  (
   );
    initial $display("%m not yet modelled!!");
endmodule // sn74ls74
