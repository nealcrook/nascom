//
module sn74ls32
  (
   output p11,
   output p8,
//   output p8,
//   output p11,

   input  p12,
   input  p13,

   input  p9,
   input  p10

//   input  p9,
//   input  p10,

//   input  p12,
//   input  p13
   );



endmodule // sn74ls32
