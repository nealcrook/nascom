//
module mk4118
  (// Input/Output
   inout d7,
   inout d6,
   inout d5,
   inout d4,
   inout d3,
   inout d2,
   inout d1,
   inout d0,
   // In
   input a9,
   input a8,
   input a7,
   input a6,
   input a5,
   input a4,
   input a3,
   input a2,
   input a1,
   input a0,
   //
   input ce_n,
   input we_n,
   input oe_n
   );

    initial $display("%m not yet modelled!!");
endmodule // mk4118



