//
module sn74ls14
  (
   );
    initial $display("%m not yet modelled!!");
endmodule // sn74ls14

