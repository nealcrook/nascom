//
module eprom2716
  (
   );
    initial $display("%m not yet modelled!!");
endmodule // eprom2716

