//
module sn81ls97
  (
   output p17,
   output p3,
   output p5,
   output p7,
   output p9,
   output p11,
   output p13,
   output p15,

   input  p18,
   input  p2,
   input  p4,
   input  p6,
   input  p8,
   input  p12,
   input  p14,
   input  p16,

   input  p1,
   input  p19
   );

endmodule // sn81ls97
