//
module mk4118
  (
   );
    initial $display("%m not yet modelled!!");
endmodule // mk4118



