//
module dp8304
  (// In/Out
   inout p8,
   inout p1,
   inout p2,
   inout p3,
   inout p4,
   inout p5,
   inout p6,
   inout p7,
   //
   inout p12,
   inout p19,
   inout p18,
   inout p17,
   inout p16,
   inout p15,
   inout p14,
   inout p13,
   // In
   input p11_dir,
   input p9_g
   );
    initial $display("%m not yet modelled!!");
endmodule // dp8304

