//
module sn74ls10
  (
   );
    initial $display("%m not yet modelled!!");
endmodule // sn74ls10
